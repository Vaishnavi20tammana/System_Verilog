class transaction;
  rand logic d;
  logic q;
  logic q_expected;
  
endclass
